`ifndef sprites_vh
`define sprites_vh

`define APPLE_PIC \
sp[0][0][0] = 3'b111;\
sp[0][0][1] = 3'b111;\
sp[0][0][2] = 3'b111;\
sp[0][0][3] = 3'b111;\
sp[0][0][4] = 3'b000;\
sp[0][0][5] = 3'b000;\
sp[0][0][6] = 3'b000;\
sp[0][0][7] = 3'b000;\
sp[0][0][8] = 3'b000;\
sp[0][0][9] = 3'b000;\
sp[0][0][10] = 3'b000;\
sp[0][0][11] = 3'b000;\
sp[0][0][12] = 3'b111;\
sp[0][0][13] = 3'b111;\
sp[0][0][14] = 3'b111;\
sp[0][0][15] = 3'b111;\
sp[0][1][0] = 3'b111;\
sp[0][1][1] = 3'b111;\
sp[0][1][2] = 3'b111;\
sp[0][1][3] = 3'b000;\
sp[0][1][4] = 3'b100;\
sp[0][1][5] = 3'b100;\
sp[0][1][6] = 3'b100;\
sp[0][1][7] = 3'b100;\
sp[0][1][8] = 3'b100;\
sp[0][1][9] = 3'b100;\
sp[0][1][10] = 3'b100;\
sp[0][1][11] = 3'b100;\
sp[0][1][12] = 3'b000;\
sp[0][1][13] = 3'b111;\
sp[0][1][14] = 3'b111;\
sp[0][1][15] = 3'b111;\
sp[0][2][0] = 3'b111;\
sp[0][2][1] = 3'b111;\
sp[0][2][2] = 3'b000;\
sp[0][2][3] = 3'b100;\
sp[0][2][4] = 3'b100;\
sp[0][2][5] = 3'b000;\
sp[0][2][6] = 3'b000;\
sp[0][2][7] = 3'b000;\
sp[0][2][8] = 3'b100;\
sp[0][2][9] = 3'b100;\
sp[0][2][10] = 3'b100;\
sp[0][2][11] = 3'b100;\
sp[0][2][12] = 3'b100;\
sp[0][2][13] = 3'b000;\
sp[0][2][14] = 3'b111;\
sp[0][2][15] = 3'b111;\
sp[0][3][0] = 3'b111;\
sp[0][3][1] = 3'b000;\
sp[0][3][2] = 3'b100;\
sp[0][3][3] = 3'b100;\
sp[0][3][4] = 3'b000;\
sp[0][3][5] = 3'b000;\
sp[0][3][6] = 3'b000;\
sp[0][3][7] = 3'b000;\
sp[0][3][8] = 3'b100;\
sp[0][3][9] = 3'b100;\
sp[0][3][10] = 3'b100;\
sp[0][3][11] = 3'b100;\
sp[0][3][12] = 3'b100;\
sp[0][3][13] = 3'b100;\
sp[0][3][14] = 3'b000;\
sp[0][3][15] = 3'b111;\
sp[0][4][0] = 3'b000;\
sp[0][4][1] = 3'b100;\
sp[0][4][2] = 3'b100;\
sp[0][4][3] = 3'b000;\
sp[0][4][4] = 3'b010;\
sp[0][4][5] = 3'b010;\
sp[0][4][6] = 3'b010;\
sp[0][4][7] = 3'b000;\
sp[0][4][8] = 3'b100;\
sp[0][4][9] = 3'b100;\
sp[0][4][10] = 3'b100;\
sp[0][4][11] = 3'b100;\
sp[0][4][12] = 3'b100;\
sp[0][4][13] = 3'b100;\
sp[0][4][14] = 3'b100;\
sp[0][4][15] = 3'b000;\
sp[0][5][0] = 3'b000;\
sp[0][5][1] = 3'b100;\
sp[0][5][2] = 3'b000;\
sp[0][5][3] = 3'b010;\
sp[0][5][4] = 3'b010;\
sp[0][5][5] = 3'b010;\
sp[0][5][6] = 3'b010;\
sp[0][5][7] = 3'b000;\
sp[0][5][8] = 3'b100;\
sp[0][5][9] = 3'b100;\
sp[0][5][10] = 3'b100;\
sp[0][5][11] = 3'b100;\
sp[0][5][12] = 3'b100;\
sp[0][5][13] = 3'b100;\
sp[0][5][14] = 3'b100;\
sp[0][5][15] = 3'b000;\
sp[0][6][0] = 3'b000;\
sp[0][6][1] = 3'b100;\
sp[0][6][2] = 3'b000;\
sp[0][6][3] = 3'b010;\
sp[0][6][4] = 3'b010;\
sp[0][6][5] = 3'b010;\
sp[0][6][6] = 3'b000;\
sp[0][6][7] = 3'b100;\
sp[0][6][8] = 3'b100;\
sp[0][6][9] = 3'b100;\
sp[0][6][10] = 3'b100;\
sp[0][6][11] = 3'b100;\
sp[0][6][12] = 3'b100;\
sp[0][6][13] = 3'b100;\
sp[0][6][14] = 3'b100;\
sp[0][6][15] = 3'b000;\
sp[0][7][0] = 3'b000;\
sp[0][7][1] = 3'b000;\
sp[0][7][2] = 3'b000;\
sp[0][7][3] = 3'b000;\
sp[0][7][4] = 3'b000;\
sp[0][7][5] = 3'b000;\
sp[0][7][6] = 3'b100;\
sp[0][7][7] = 3'b100;\
sp[0][7][8] = 3'b100;\
sp[0][7][9] = 3'b100;\
sp[0][7][10] = 3'b100;\
sp[0][7][11] = 3'b100;\
sp[0][7][12] = 3'b100;\
sp[0][7][13] = 3'b100;\
sp[0][7][14] = 3'b100;\
sp[0][7][15] = 3'b000;\
sp[0][8][0] = 3'b000;\
sp[0][8][1] = 3'b000;\
sp[0][8][2] = 3'b000;\
sp[0][8][3] = 3'b100;\
sp[0][8][4] = 3'b100;\
sp[0][8][5] = 3'b100;\
sp[0][8][6] = 3'b100;\
sp[0][8][7] = 3'b100;\
sp[0][8][8] = 3'b100;\
sp[0][8][9] = 3'b100;\
sp[0][8][10] = 3'b100;\
sp[0][8][11] = 3'b100;\
sp[0][8][12] = 3'b100;\
sp[0][8][13] = 3'b100;\
sp[0][8][14] = 3'b100;\
sp[0][8][15] = 3'b000;\
sp[0][9][0] = 3'b000;\
sp[0][9][1] = 3'b100;\
sp[0][9][2] = 3'b100;\
sp[0][9][3] = 3'b100;\
sp[0][9][4] = 3'b100;\
sp[0][9][5] = 3'b100;\
sp[0][9][6] = 3'b100;\
sp[0][9][7] = 3'b100;\
sp[0][9][8] = 3'b100;\
sp[0][9][9] = 3'b100;\
sp[0][9][10] = 3'b100;\
sp[0][9][11] = 3'b100;\
sp[0][9][12] = 3'b100;\
sp[0][9][13] = 3'b100;\
sp[0][9][14] = 3'b100;\
sp[0][9][15] = 3'b000;\
sp[0][10][0] = 3'b000;\
sp[0][10][1] = 3'b100;\
sp[0][10][2] = 3'b100;\
sp[0][10][3] = 3'b100;\
sp[0][10][4] = 3'b100;\
sp[0][10][5] = 3'b100;\
sp[0][10][6] = 3'b111;\
sp[0][10][7] = 3'b111;\
sp[0][10][8] = 3'b111;\
sp[0][10][9] = 3'b100;\
sp[0][10][10] = 3'b100;\
sp[0][10][11] = 3'b100;\
sp[0][10][12] = 3'b100;\
sp[0][10][13] = 3'b100;\
sp[0][10][14] = 3'b100;\
sp[0][10][15] = 3'b000;\
sp[0][11][0] = 3'b000;\
sp[0][11][1] = 3'b100;\
sp[0][11][2] = 3'b100;\
sp[0][11][3] = 3'b100;\
sp[0][11][4] = 3'b100;\
sp[0][11][5] = 3'b111;\
sp[0][11][6] = 3'b111;\
sp[0][11][7] = 3'b111;\
sp[0][11][8] = 3'b111;\
sp[0][11][9] = 3'b111;\
sp[0][11][10] = 3'b100;\
sp[0][11][11] = 3'b100;\
sp[0][11][12] = 3'b100;\
sp[0][11][13] = 3'b100;\
sp[0][11][14] = 3'b100;\
sp[0][11][15] = 3'b000;\
sp[0][12][0] = 3'b000;\
sp[0][12][1] = 3'b100;\
sp[0][12][2] = 3'b100;\
sp[0][12][3] = 3'b100;\
sp[0][12][4] = 3'b100;\
sp[0][12][5] = 3'b100;\
sp[0][12][6] = 3'b111;\
sp[0][12][7] = 3'b111;\
sp[0][12][8] = 3'b111;\
sp[0][12][9] = 3'b100;\
sp[0][12][10] = 3'b100;\
sp[0][12][11] = 3'b100;\
sp[0][12][12] = 3'b100;\
sp[0][12][13] = 3'b100;\
sp[0][12][14] = 3'b100;\
sp[0][12][15] = 3'b000;\
sp[0][13][0] = 3'b111;\
sp[0][13][1] = 3'b111;\
sp[0][13][2] = 3'b000;\
sp[0][13][3] = 3'b100;\
sp[0][13][4] = 3'b100;\
sp[0][13][5] = 3'b100;\
sp[0][13][6] = 3'b100;\
sp[0][13][7] = 3'b100;\
sp[0][13][8] = 3'b100;\
sp[0][13][9] = 3'b100;\
sp[0][13][10] = 3'b100;\
sp[0][13][11] = 3'b100;\
sp[0][13][12] = 3'b100;\
sp[0][13][13] = 3'b000;\
sp[0][13][14] = 3'b111;\
sp[0][13][15] = 3'b111;\
sp[0][14][0] = 3'b111;\
sp[0][14][1] = 3'b111;\
sp[0][14][2] = 3'b111;\
sp[0][14][3] = 3'b000;\
sp[0][14][4] = 3'b100;\
sp[0][14][5] = 3'b100;\
sp[0][14][6] = 3'b100;\
sp[0][14][7] = 3'b100;\
sp[0][14][8] = 3'b100;\
sp[0][14][9] = 3'b100;\
sp[0][14][10] = 3'b100;\
sp[0][14][11] = 3'b100;\
sp[0][14][12] = 3'b000;\
sp[0][14][13] = 3'b111;\
sp[0][14][14] = 3'b111;\
sp[0][14][15] = 3'b111;\
sp[0][15][0] = 3'b111;\
sp[0][15][1] = 3'b111;\
sp[0][15][2] = 3'b111;\
sp[0][15][3] = 3'b111;\
sp[0][15][4] = 3'b000;\
sp[0][15][5] = 3'b000;\
sp[0][15][6] = 3'b000;\
sp[0][15][7] = 3'b000;\
sp[0][15][8] = 3'b000;\
sp[0][15][9] = 3'b000;\
sp[0][15][10] = 3'b000;\
sp[0][15][11] = 3'b000;\
sp[0][15][12] = 3'b111;\
sp[0][15][13] = 3'b111;\
sp[0][15][14] = 3'b111;\
sp[0][15][15] = 3'b111;\
`define SPRITE_INIT `APPLE_PIC

`endif // sprites_vh