define Gift 
sp[0][0][0] = 3'b000;\
sp[0][0][1] = 3'b000;\
sp[0][0][2] = 3'b000;\
sp[0][0][3] = 3'b000;\
sp[0][0][4] = 3'b000;\
sp[0][0][5] = 3'b000;\
sp[0][0][6] = 3'b000;\
sp[0][0][7] = 3'b000;\
sp[0][0][8] = 3'b000;\
sp[0][0][9] = 3'b000;\
sp[0][0][10] = 3'b000;\
sp[0][0][11] = 3'b000;\
sp[0][0][12] = 3'b000;\
sp[0][0][13] = 3'b000;\
sp[0][0][14] = 3'b000;\
sp[0][0][15] = 3'b000;\
sp[0][1][0] = 3'b000;\
sp[0][1][1] = 3'b100;\
sp[0][1][2] = 3'b100;\
sp[0][1][3] = 3'b100;\
sp[0][1][4] = 3'b100;\
sp[0][1][5] = 3'b100;\
sp[0][1][6] = 3'b100;\
sp[0][1][7] = 3'b111;\
sp[0][1][8] = 3'b111;\
sp[0][1][9] = 3'b100;\
sp[0][1][10] = 3'b100;\
sp[0][1][11] = 3'b100;\
sp[0][1][12] = 3'b100;\
sp[0][1][13] = 3'b100;\
sp[0][1][14] = 3'b100;\
sp[0][1][15] = 3'b000;\
sp[0][2][0] = 3'b000;\
sp[0][2][1] = 3'b100;\
sp[0][2][2] = 3'b100;\
sp[0][2][3] = 3'b100;\
sp[0][2][4] = 3'b100;\
sp[0][2][5] = 3'b100;\
sp[0][2][6] = 3'b100;\
sp[0][2][7] = 3'b111;\
sp[0][2][8] = 3'b111;\
sp[0][2][9] = 3'b100;\
sp[0][2][10] = 3'b100;\
sp[0][2][11] = 3'b100;\
sp[0][2][12] = 3'b100;\
sp[0][2][13] = 3'b100;\
sp[0][2][14] = 3'b100;\
sp[0][2][15] = 3'b000;\
sp[0][3][0] = 3'b000;\
sp[0][3][1] = 3'b100;\
sp[0][3][2] = 3'b100;\
sp[0][3][3] = 3'b100;\
sp[0][3][4] = 3'b100;\
sp[0][3][5] = 3'b100;\
sp[0][3][6] = 3'b100;\
sp[0][3][7] = 3'b111;\
sp[0][3][8] = 3'b111;\
sp[0][3][9] = 3'b100;\
sp[0][3][10] = 3'b100;\
sp[0][3][11] = 3'b100;\
sp[0][3][12] = 3'b100;\
sp[0][3][13] = 3'b100;\
sp[0][3][14] = 3'b100;\
sp[0][3][15] = 3'b000;\
sp[0][4][0] = 3'b000;\
sp[0][4][1] = 3'b100;\
sp[0][4][2] = 3'b100;\
sp[0][4][3] = 3'b100;\
sp[0][4][4] = 3'b100;\
sp[0][4][5] = 3'b100;\
sp[0][4][6] = 3'b100;\
sp[0][4][7] = 3'b111;\
sp[0][4][8] = 3'b111;\
sp[0][4][9] = 3'b100;\
sp[0][4][10] = 3'b100;\
sp[0][4][11] = 3'b100;\
sp[0][4][12] = 3'b100;\
sp[0][4][13] = 3'b100;\
sp[0][4][14] = 3'b100;\
sp[0][4][15] = 3'b000;\
sp[0][5][0] = 3'b000;\
sp[0][5][1] = 3'b100;\
sp[0][5][2] = 3'b100;\
sp[0][5][3] = 3'b100;\
sp[0][5][4] = 3'b100;\
sp[0][5][5] = 3'b100;\
sp[0][5][6] = 3'b100;\
sp[0][5][7] = 3'b111;\
sp[0][5][8] = 3'b111;\
sp[0][5][9] = 3'b100;\
sp[0][5][10] = 3'b100;\
sp[0][5][11] = 3'b100;\
sp[0][5][12] = 3'b100;\
sp[0][5][13] = 3'b100;\
sp[0][5][14] = 3'b100;\
sp[0][5][15] = 3'b000;\
sp[0][6][0] = 3'b000;\
sp[0][6][1] = 3'b100;\
sp[0][6][2] = 3'b100;\
sp[0][6][3] = 3'b100;\
sp[0][6][4] = 3'b100;\
sp[0][6][5] = 3'b100;\
sp[0][6][6] = 3'b100;\
sp[0][6][7] = 3'b111;\
sp[0][6][8] = 3'b111;\
sp[0][6][9] = 3'b100;\
sp[0][6][10] = 3'b100;\
sp[0][6][11] = 3'b100;\
sp[0][6][12] = 3'b100;\
sp[0][6][13] = 3'b100;\
sp[0][6][14] = 3'b100;\
sp[0][6][15] = 3'b000;\
sp[0][7][0] = 3'b000;\
sp[0][7][1] = 3'b111;\
sp[0][7][2] = 3'b111;\
sp[0][7][3] = 3'b111;\
sp[0][7][4] = 3'b111;\
sp[0][7][5] = 3'b111;\
sp[0][7][6] = 3'b111;\
sp[0][7][7] = 3'b111;\
sp[0][7][8] = 3'b111;\
sp[0][7][9] = 3'b111;\
sp[0][7][10] = 3'b111;\
sp[0][7][11] = 3'b111;\
sp[0][7][12] = 3'b111;\
sp[0][7][13] = 3'b111;\
sp[0][7][14] = 3'b111;\
sp[0][7][15] = 3'b000;\
sp[0][8][0] = 3'b000;\
sp[0][8][1] = 3'b111;\
sp[0][8][2] = 3'b111;\
sp[0][8][3] = 3'b111;\
sp[0][8][4] = 3'b111;\
sp[0][8][5] = 3'b111;\
sp[0][8][6] = 3'b111;\
sp[0][8][7] = 3'b111;\
sp[0][8][8] = 3'b111;\
sp[0][8][9] = 3'b111;\
sp[0][8][10] = 3'b111;\
sp[0][8][11] = 3'b111;\
sp[0][8][12] = 3'b111;\
sp[0][8][13] = 3'b111;\
sp[0][8][14] = 3'b111;\
sp[0][8][15] = 3'b000;\
sp[0][9][0] = 3'b000;\
sp[0][9][1] = 3'b100;\
sp[0][9][2] = 3'b100;\
sp[0][9][3] = 3'b100;\
sp[0][9][4] = 3'b100;\
sp[0][9][5] = 3'b100;\
sp[0][9][6] = 3'b100;\
sp[0][9][7] = 3'b111;\
sp[0][9][8] = 3'b111;\
sp[0][9][9] = 3'b100;\
sp[0][9][10] = 3'b100;\
sp[0][9][11] = 3'b100;\
sp[0][9][12] = 3'b100;\
sp[0][9][13] = 3'b100;\
sp[0][9][14] = 3'b100;\
sp[0][9][15] = 3'b000;\
sp[0][10][0] = 3'b000;\
sp[0][10][1] = 3'b100;\
sp[0][10][2] = 3'b100;\
sp[0][10][3] = 3'b100;\
sp[0][10][4] = 3'b100;\
sp[0][10][5] = 3'b100;\
sp[0][10][6] = 3'b100;\
sp[0][10][7] = 3'b111;\
sp[0][10][8] = 3'b111;\
sp[0][10][9] = 3'b100;\
sp[0][10][10] = 3'b100;\
sp[0][10][11] = 3'b100;\
sp[0][10][12] = 3'b100;\
sp[0][10][13] = 3'b100;\
sp[0][10][14] = 3'b100;\
sp[0][10][15] = 3'b000;\
sp[0][11][0] = 3'b000;\
sp[0][11][1] = 3'b100;\
sp[0][11][2] = 3'b100;\
sp[0][11][3] = 3'b100;\
sp[0][11][4] = 3'b100;\
sp[0][11][5] = 3'b100;\
sp[0][11][6] = 3'b100;\
sp[0][11][7] = 3'b111;\
sp[0][11][8] = 3'b111;\
sp[0][11][9] = 3'b100;\
sp[0][11][10] = 3'b100;\
sp[0][11][11] = 3'b100;\
sp[0][11][12] = 3'b100;\
sp[0][11][13] = 3'b100;\
sp[0][11][14] = 3'b100;\
sp[0][11][15] = 3'b000;\
sp[0][12][0] = 3'b000;\
sp[0][12][1] = 3'b100;\
sp[0][12][2] = 3'b100;\
sp[0][12][3] = 3'b100;\
sp[0][12][4] = 3'b100;\
sp[0][12][5] = 3'b100;\
sp[0][12][6] = 3'b100;\
sp[0][12][7] = 3'b111;\
sp[0][12][8] = 3'b111;\
sp[0][12][9] = 3'b100;\
sp[0][12][10] = 3'b100;\
sp[0][12][11] = 3'b100;\
sp[0][12][12] = 3'b100;\
sp[0][12][13] = 3'b100;\
sp[0][12][14] = 3'b100;\
sp[0][12][15] = 3'b000;\
sp[0][13][0] = 3'b000;\
sp[0][13][1] = 3'b100;\
sp[0][13][2] = 3'b100;\
sp[0][13][3] = 3'b100;\
sp[0][13][4] = 3'b100;\
sp[0][13][5] = 3'b100;\
sp[0][13][6] = 3'b100;\
sp[0][13][7] = 3'b111;\
sp[0][13][8] = 3'b111;\
sp[0][13][9] = 3'b100;\
sp[0][13][10] = 3'b100;\
sp[0][13][11] = 3'b100;\
sp[0][13][12] = 3'b100;\
sp[0][13][13] = 3'b100;\
sp[0][13][14] = 3'b100;\
sp[0][13][15] = 3'b000;\
sp[0][14][0] = 3'b000;\
sp[0][14][1] = 3'b100;\
sp[0][14][2] = 3'b100;\
sp[0][14][3] = 3'b100;\
sp[0][14][4] = 3'b100;\
sp[0][14][5] = 3'b100;\
sp[0][14][6] = 3'b100;\
sp[0][14][7] = 3'b111;\
sp[0][14][8] = 3'b111;\
sp[0][14][9] = 3'b100;\
sp[0][14][10] = 3'b100;\
sp[0][14][11] = 3'b100;\
sp[0][14][12] = 3'b100;\
sp[0][14][13] = 3'b100;\
sp[0][14][14] = 3'b100;\
sp[0][14][15] = 3'b000;\
sp[0][15][0] = 3'b000;\
sp[0][15][1] = 3'b000;\
sp[0][15][2] = 3'b000;\
sp[0][15][3] = 3'b000;\
sp[0][15][4] = 3'b000;\
sp[0][15][5] = 3'b000;\
sp[0][15][6] = 3'b000;\
sp[0][15][7] = 3'b000;\
sp[0][15][8] = 3'b000;\
sp[0][15][9] = 3'b000;\
sp[0][15][10] = 3'b000;\
sp[0][15][11] = 3'b000;\
sp[0][15][12] = 3'b000;\
sp[0][15][13] = 3'b000;\
sp[0][15][14] = 3'b000;\
sp[0][15][15] = 3'b000;\
define Grinch \
sp[1][0][0] = 3'b111;\
sp[1][0][1] = 3'b111;\
sp[1][0][2] = 3'b111;\
sp[1][0][3] = 3'b111;\
sp[1][0][4] = 3'b111;\
sp[1][0][5] = 3'b111;\
sp[1][0][6] = 3'b111;\
sp[1][0][7] = 3'b111;\
sp[1][0][8] = 3'b111;\
sp[1][0][9] = 3'b111;\
sp[1][0][10] = 3'b111;\
sp[1][0][11] = 3'b111;\
sp[1][0][12] = 3'b111;\
sp[1][0][13] = 3'b111;\
sp[1][0][14] = 3'b111;\
sp[1][0][15] = 3'b111;\
sp[1][1][0] = 3'b111;\
sp[1][1][1] = 3'b111;\
sp[1][1][2] = 3'b111;\
sp[1][1][3] = 3'b111;\
sp[1][1][4] = 3'b111;\
sp[1][1][5] = 3'b111;\
sp[1][1][6] = 3'b111;\
sp[1][1][7] = 3'b111;\
sp[1][1][8] = 3'b111;\
sp[1][1][9] = 3'b111;\
sp[1][1][10] = 3'b111;\
sp[1][1][11] = 3'b111;\
sp[1][1][12] = 3'b111;\
sp[1][1][13] = 3'b111;\
sp[1][1][14] = 3'b111;\
sp[1][1][15] = 3'b111;\
sp[1][2][0] = 3'b111;\
sp[1][2][1] = 3'b111;\
sp[1][2][2] = 3'b111;\
sp[1][2][3] = 3'b111;\
sp[1][2][4] = 3'b111;\
sp[1][2][5] = 3'b111;\
sp[1][2][6] = 3'b111;\
sp[1][2][7] = 3'b111;\
sp[1][2][8] = 3'b111;\
sp[1][2][9] = 3'b000;\
sp[1][2][10] = 3'b000;\
sp[1][2][11] = 3'b000;\
sp[1][2][12] = 3'b111;\
sp[1][2][13] = 3'b111;\
sp[1][2][14] = 3'b111;\
sp[1][2][15] = 3'b111;\
sp[1][3][0] = 3'b111;\
sp[1][3][1] = 3'b111;\
sp[1][3][2] = 3'b111;\
sp[1][3][3] = 3'b111;\
sp[1][3][4] = 3'b111;\
sp[1][3][5] = 3'b000;\
sp[1][3][6] = 3'b000;\
sp[1][3][7] = 3'b000;\
sp[1][3][8] = 3'b000;\
sp[1][3][9] = 3'b010;\
sp[1][3][10] = 3'b000;\
sp[1][3][11] = 3'b010;\
sp[1][3][12] = 3'b000;\
sp[1][3][13] = 3'b111;\
sp[1][3][14] = 3'b000;\
sp[1][3][15] = 3'b111;\
sp[1][4][0] = 3'b111;\
sp[1][4][1] = 3'b111;\
sp[1][4][2] = 3'b111;\
sp[1][4][3] = 3'b111;\
sp[1][4][4] = 3'b000;\
sp[1][4][5] = 3'b010;\
sp[1][4][6] = 3'b010;\
sp[1][4][7] = 3'b010;\
sp[1][4][8] = 3'b010;\
sp[1][4][9] = 3'b000;\
sp[1][4][10] = 3'b010;\
sp[1][4][11] = 3'b000;\
sp[1][4][12] = 3'b010;\
sp[1][4][13] = 3'b000;\
sp[1][4][14] = 3'b111;\
sp[1][4][15] = 3'b111;\
sp[1][5][0] = 3'b111;\
sp[1][5][1] = 3'b111;\
sp[1][5][2] = 3'b000;\
sp[1][5][3] = 3'b000;\
sp[1][5][4] = 3'b010;\
sp[1][5][5] = 3'b000;\
sp[1][5][6] = 3'b111;\
sp[1][5][7] = 3'b111;\
sp[1][5][8] = 3'b000;\
sp[1][5][9] = 3'b010;\
sp[1][5][10] = 3'b000;\
sp[1][5][11] = 3'b010;\
sp[1][5][12] = 3'b000;\
sp[1][5][13] = 3'b000;\
sp[1][5][14] = 3'b000;\
sp[1][5][15] = 3'b000;\
sp[1][6][0] = 3'b000;\
sp[1][6][1] = 3'b000;\
sp[1][6][2] = 3'b000;\
sp[1][6][3] = 3'b010;\
sp[1][6][4] = 3'b000;\
sp[1][6][5] = 3'b010;\
sp[1][6][6] = 3'b000;\
sp[1][6][7] = 3'b111;\
sp[1][6][8] = 3'b010;\
sp[1][6][9] = 3'b000;\
sp[1][6][10] = 3'b010;\
sp[1][6][11] = 3'b000;\
sp[1][6][12] = 3'b010;\
sp[1][6][13] = 3'b010;\
sp[1][6][14] = 3'b000;\
sp[1][6][15] = 3'b000;\
sp[1][7][0] = 3'b000;\
sp[1][7][1] = 3'b100;\
sp[1][7][2] = 3'b010;\
sp[1][7][3] = 3'b000;\
sp[1][7][4] = 3'b010;\
sp[1][7][5] = 3'b000;\
sp[1][7][6] = 3'b010;\
sp[1][7][7] = 3'b000;\
sp[1][7][8] = 3'b000;\
sp[1][7][9] = 3'b010;\
sp[1][7][10] = 3'b000;\
sp[1][7][11] = 3'b010;\
sp[1][7][12] = 3'b000;\
sp[1][7][13] = 3'b010;\
sp[1][7][14] = 3'b010;\
sp[1][7][15] = 3'b000;\
sp[1][8][0] = 3'b000;\
sp[1][8][1] = 3'b100;\
sp[1][8][2] = 3'b010;\
sp[1][8][3] = 3'b000;\
sp[1][8][4] = 3'b010;\
sp[1][8][5] = 3'b000;\
sp[1][8][6] = 3'b010;\
sp[1][8][7] = 3'b000;\
sp[1][8][8] = 3'b000;\
sp[1][8][9] = 3'b010;\
sp[1][8][10] = 3'b000;\
sp[1][8][11] = 3'b010;\
sp[1][8][12] = 3'b000;\
sp[1][8][13] = 3'b010;\
sp[1][8][14] = 3'b010;\
sp[1][8][15] = 3'b000;\
sp[1][9][0] = 3'b000;\
sp[1][9][1] = 3'b000;\
sp[1][9][2] = 3'b000;\
sp[1][9][3] = 3'b010;\
sp[1][9][4] = 3'b000;\
sp[1][9][5] = 3'b010;\
sp[1][9][6] = 3'b000;\
sp[1][9][7] = 3'b111;\
sp[1][9][8] = 3'b010;\
sp[1][9][9] = 3'b000;\
sp[1][9][10] = 3'b010;\
sp[1][9][11] = 3'b000;\
sp[1][9][12] = 3'b010;\
sp[1][9][13] = 3'b010;\
sp[1][9][14] = 3'b000;\
sp[1][9][15] = 3'b000;\
sp[1][10][0] = 3'b111;\
sp[1][10][1] = 3'b111;\
sp[1][10][2] = 3'b000;\
sp[1][10][3] = 3'b000;\
sp[1][10][4] = 3'b010;\
sp[1][10][5] = 3'b000;\
sp[1][10][6] = 3'b111;\
sp[1][10][7] = 3'b111;\
sp[1][10][8] = 3'b000;\
sp[1][10][9] = 3'b010;\
sp[1][10][10] = 3'b000;\
sp[1][10][11] = 3'b010;\
sp[1][10][12] = 3'b000;\
sp[1][10][13] = 3'b000;\
sp[1][10][14] = 3'b000;\
sp[1][10][15] = 3'b000;\
sp[1][11][0] = 3'b111;\
sp[1][11][1] = 3'b111;\
sp[1][11][2] = 3'b111;\
sp[1][11][3] = 3'b111;\
sp[1][11][4] = 3'b000;\
sp[1][11][5] = 3'b010;\
sp[1][11][6] = 3'b010;\
sp[1][11][7] = 3'b010;\
sp[1][11][8] = 3'b010;\
sp[1][11][9] = 3'b000;\
sp[1][11][10] = 3'b010;\
sp[1][11][11] = 3'b000;\
sp[1][11][12] = 3'b010;\
sp[1][11][13] = 3'b000;\
sp[1][11][14] = 3'b111;\
sp[1][11][15] = 3'b111;\
sp[1][12][0] = 3'b111;\
sp[1][12][1] = 3'b111;\
sp[1][12][2] = 3'b111;\
sp[1][12][3] = 3'b111;\
sp[1][12][4] = 3'b111;\
sp[1][12][5] = 3'b000;\
sp[1][12][6] = 3'b000;\
sp[1][12][7] = 3'b000;\
sp[1][12][8] = 3'b000;\
sp[1][12][9] = 3'b010;\
sp[1][12][10] = 3'b000;\
sp[1][12][11] = 3'b010;\
sp[1][12][12] = 3'b000;\
sp[1][12][13] = 3'b111;\
sp[1][12][14] = 3'b000;\
sp[1][12][15] = 3'b111;\
sp[1][13][0] = 3'b111;\
sp[1][13][1] = 3'b111;\
sp[1][13][2] = 3'b111;\
sp[1][13][3] = 3'b111;\
sp[1][13][4] = 3'b111;\
sp[1][13][5] = 3'b111;\
sp[1][13][6] = 3'b111;\
sp[1][13][7] = 3'b111;\
sp[1][13][8] = 3'b111;\
sp[1][13][9] = 3'b000;\
sp[1][13][10] = 3'b000;\
sp[1][13][11] = 3'b000;\
sp[1][13][12] = 3'b111;\
sp[1][13][13] = 3'b111;\
sp[1][13][14] = 3'b111;\
sp[1][13][15] = 3'b111;\
sp[1][14][0] = 3'b111;\
sp[1][14][1] = 3'b111;\
sp[1][14][2] = 3'b111;\
sp[1][14][3] = 3'b111;\
sp[1][14][4] = 3'b111;\
sp[1][14][5] = 3'b111;\
sp[1][14][6] = 3'b111;\
sp[1][14][7] = 3'b111;\
sp[1][14][8] = 3'b111;\
sp[1][14][9] = 3'b111;\
sp[1][14][10] = 3'b111;\
sp[1][14][11] = 3'b111;\
sp[1][14][12] = 3'b111;\
sp[1][14][13] = 3'b111;\
sp[1][14][14] = 3'b111;\
sp[1][14][15] = 3'b111;\
sp[1][15][0] = 3'b111;\
sp[1][15][1] = 3'b111;\
sp[1][15][2] = 3'b111;\
sp[1][15][3] = 3'b111;\
sp[1][15][4] = 3'b111;\
sp[1][15][5] = 3'b111;\
sp[1][15][6] = 3'b111;\
sp[1][15][7] = 3'b111;\
sp[1][15][8] = 3'b111;\
sp[1][15][9] = 3'b111;\
sp[1][15][10] = 3'b111;\
sp[1][15][11] = 3'b111;\
sp[1][15][12] = 3'b111;\
sp[1][15][13] = 3'b111;\
sp[1][15][14] = 3'b111;\
sp[1][15][15] = 3'b111;\

/////Wall
sp[2][0][0] = 3'b000;\
sp[2][0][1] = 3'b000;\
sp[2][0][2] = 3'b000;\
sp[2][0][3] = 3'b111;\
sp[2][0][4] = 3'b111;\
sp[2][0][5] = 3'b000;\
sp[2][0][6] = 3'b000;\
sp[2][0][7] = 3'b000;\
sp[2][0][8] = 3'b000;\
sp[2][0][9] = 3'b111;\
sp[2][0][10] = 3'b111;\
sp[2][0][11] = 3'b000;\
sp[2][0][12] = 3'b000;\
sp[2][0][13] = 3'b000;\
sp[2][0][14] = 3'b000;\
sp[2][0][15] = 3'b000;\
sp[2][1][0] = 3'b000;\
sp[2][1][1] = 3'b111;\
sp[2][1][2] = 3'b111;\
sp[2][1][3] = 3'b000;\
sp[2][1][4] = 3'b000;\
sp[2][1][5] = 3'b111;\
sp[2][1][6] = 3'b111;\
sp[2][1][7] = 3'b000;\
sp[2][1][8] = 3'b000;\
sp[2][1][9] = 3'b111;\
sp[2][1][10] = 3'b111;\
sp[2][1][11] = 3'b000;\
sp[2][1][12] = 3'b111;\
sp[2][1][13] = 3'b111;\
sp[2][1][14] = 3'b000;\
sp[2][1][15] = 3'b000;\
sp[2][2][0] = 3'b000;\
sp[2][2][1] = 3'b111;\
sp[2][2][2] = 3'b111;\
sp[2][2][3] = 3'b000;\
sp[2][2][4] = 3'b000;\
sp[2][2][5] = 3'b111;\
sp[2][2][6] = 3'b111;\
sp[2][2][7] = 3'b000;\
sp[2][2][8] = 3'b000;\
sp[2][2][9] = 3'b111;\
sp[2][2][10] = 3'b111;\
sp[2][2][11] = 3'b000;\
sp[2][2][12] = 3'b111;\
sp[2][2][13] = 3'b111;\
sp[2][2][14] = 3'b000;\
sp[2][2][15] = 3'b000;\
sp[2][3][0] = 3'b000;\
sp[2][3][1] = 3'b000;\
sp[2][3][2] = 3'b000;\
sp[2][3][3] = 3'b111;\
sp[2][3][4] = 3'b111;\
sp[2][3][5] = 3'b000;\
sp[2][3][6] = 3'b000;\
sp[2][3][7] = 3'b000;\
sp[2][3][8] = 3'b000;\
sp[2][3][9] = 3'b111;\
sp[2][3][10] = 3'b111;\
sp[2][3][11] = 3'b000;\
sp[2][3][12] = 3'b000;\
sp[2][3][13] = 3'b000;\
sp[2][3][14] = 3'b000;\
sp[2][3][15] = 3'b000;\
sp[2][4][0] = 3'b000;\
sp[2][4][1] = 3'b000;\
sp[2][4][2] = 3'b000;\
sp[2][4][3] = 3'b111;\
sp[2][4][4] = 3'b111;\
sp[2][4][5] = 3'b000;\
sp[2][4][6] = 3'b000;\
sp[2][4][7] = 3'b000;\
sp[2][4][8] = 3'b000;\
sp[2][4][9] = 3'b111;\
sp[2][4][10] = 3'b111;\
sp[2][4][11] = 3'b000;\
sp[2][4][12] = 3'b000;\
sp[2][4][13] = 3'b000;\
sp[2][4][14] = 3'b000;\
sp[2][4][15] = 3'b000;\
sp[2][5][0] = 3'b000;\
sp[2][5][1] = 3'b111;\
sp[2][5][2] = 3'b111;\
sp[2][5][3] = 3'b000;\
sp[2][5][4] = 3'b000;\
sp[2][5][5] = 3'b111;\
sp[2][5][6] = 3'b111;\
sp[2][5][7] = 3'b000;\
sp[2][5][8] = 3'b000;\
sp[2][5][9] = 3'b111;\
sp[2][5][10] = 3'b111;\
sp[2][5][11] = 3'b000;\
sp[2][5][12] = 3'b111;\
sp[2][5][13] = 3'b111;\
sp[2][5][14] = 3'b000;\
sp[2][5][15] = 3'b000;\
sp[2][6][0] = 3'b000;\
sp[2][6][1] = 3'b111;\
sp[2][6][2] = 3'b111;\
sp[2][6][3] = 3'b000;\
sp[2][6][4] = 3'b000;\
sp[2][6][5] = 3'b111;\
sp[2][6][6] = 3'b111;\
sp[2][6][7] = 3'b000;\
sp[2][6][8] = 3'b000;\
sp[2][6][9] = 3'b111;\
sp[2][6][10] = 3'b111;\
sp[2][6][11] = 3'b000;\
sp[2][6][12] = 3'b111;\
sp[2][6][13] = 3'b111;\
sp[2][6][14] = 3'b000;\
sp[2][6][15] = 3'b000;\
sp[2][7][0] = 3'b000;\
sp[2][7][1] = 3'b000;\
sp[2][7][2] = 3'b000;\
sp[2][7][3] = 3'b111;\
sp[2][7][4] = 3'b111;\
sp[2][7][5] = 3'b000;\
sp[2][7][6] = 3'b000;\
sp[2][7][7] = 3'b000;\
sp[2][7][8] = 3'b000;\
sp[2][7][9] = 3'b111;\
sp[2][7][10] = 3'b111;\
sp[2][7][11] = 3'b000;\
sp[2][7][12] = 3'b000;\
sp[2][7][13] = 3'b000;\
sp[2][7][14] = 3'b000;\
sp[2][7][15] = 3'b000;\
sp[2][8][0] = 3'b000;\
sp[2][8][1] = 3'b000;\
sp[2][8][2] = 3'b000;\
sp[2][8][3] = 3'b111;\
sp[2][8][4] = 3'b111;\
sp[2][8][5] = 3'b000;\
sp[2][8][6] = 3'b000;\
sp[2][8][7] = 3'b000;\
sp[2][8][8] = 3'b000;\
sp[2][8][9] = 3'b111;\
sp[2][8][10] = 3'b111;\
sp[2][8][11] = 3'b000;\
sp[2][8][12] = 3'b000;\
sp[2][8][13] = 3'b000;\
sp[2][8][14] = 3'b000;\
sp[2][8][15] = 3'b000;\
sp[2][9][0] = 3'b000;\
sp[2][9][1] = 3'b111;\
sp[2][9][2] = 3'b111;\
sp[2][9][3] = 3'b000;\
sp[2][9][4] = 3'b000;\
sp[2][9][5] = 3'b111;\
sp[2][9][6] = 3'b111;\
sp[2][9][7] = 3'b000;\
sp[2][9][8] = 3'b000;\
sp[2][9][9] = 3'b111;\
sp[2][9][10] = 3'b111;\
sp[2][9][11] = 3'b000;\
sp[2][9][12] = 3'b111;\
sp[2][9][13] = 3'b111;\
sp[2][9][14] = 3'b000;\
sp[2][9][15] = 3'b000;\
sp[2][10][0] = 3'b000;\
sp[2][10][1] = 3'b111;\
sp[2][10][2] = 3'b111;\
sp[2][10][3] = 3'b000;\
sp[2][10][4] = 3'b000;\
sp[2][10][5] = 3'b111;\
sp[2][10][6] = 3'b111;\
sp[2][10][7] = 3'b000;\
sp[2][10][8] = 3'b000;\
sp[2][10][9] = 3'b111;\
sp[2][10][10] = 3'b111;\
sp[2][10][11] = 3'b000;\
sp[2][10][12] = 3'b111;\
sp[2][10][13] = 3'b111;\
sp[2][10][14] = 3'b000;\
sp[2][10][15] = 3'b000;\
sp[2][11][0] = 3'b000;\
sp[2][11][1] = 3'b000;\
sp[2][11][2] = 3'b000;\
sp[2][11][3] = 3'b111;\
sp[2][11][4] = 3'b111;\
sp[2][11][5] = 3'b000;\
sp[2][11][6] = 3'b000;\
sp[2][11][7] = 3'b000;\
sp[2][11][8] = 3'b000;\
sp[2][11][9] = 3'b111;\
sp[2][11][10] = 3'b111;\
sp[2][11][11] = 3'b000;\
sp[2][11][12] = 3'b000;\
sp[2][11][13] = 3'b000;\
sp[2][11][14] = 3'b000;\
sp[2][11][15] = 3'b000;\
sp[2][12][0] = 3'b000;\
sp[2][12][1] = 3'b000;\
sp[2][12][2] = 3'b000;\
sp[2][12][3] = 3'b111;\
sp[2][12][4] = 3'b111;\
sp[2][12][5] = 3'b000;\
sp[2][12][6] = 3'b000;\
sp[2][12][7] = 3'b000;\
sp[2][12][8] = 3'b000;\
sp[2][12][9] = 3'b111;\
sp[2][12][10] = 3'b111;\
sp[2][12][11] = 3'b000;\
sp[2][12][12] = 3'b000;\
sp[2][12][13] = 3'b000;\
sp[2][12][14] = 3'b000;\
sp[2][12][15] = 3'b000;\
sp[2][13][0] = 3'b000;\
sp[2][13][1] = 3'b111;\
sp[2][13][2] = 3'b111;\
sp[2][13][3] = 3'b000;\
sp[2][13][4] = 3'b000;\
sp[2][13][5] = 3'b111;\
sp[2][13][6] = 3'b111;\
sp[2][13][7] = 3'b000;\
sp[2][13][8] = 3'b000;\
sp[2][13][9] = 3'b111;\
sp[2][13][10] = 3'b111;\
sp[2][13][11] = 3'b000;\
sp[2][13][12] = 3'b111;\
sp[2][13][13] = 3'b111;\
sp[2][13][14] = 3'b000;\
sp[2][13][15] = 3'b000;\
sp[2][14][0] = 3'b000;\
sp[2][14][1] = 3'b111;\
sp[2][14][2] = 3'b111;\
sp[2][14][3] = 3'b000;\
sp[2][14][4] = 3'b000;\
sp[2][14][5] = 3'b111;\
sp[2][14][6] = 3'b111;\
sp[2][14][7] = 3'b000;\
sp[2][14][8] = 3'b000;\
sp[2][14][9] = 3'b111;\
sp[2][14][10] = 3'b111;\
sp[2][14][11] = 3'b000;\
sp[2][14][12] = 3'b111;\
sp[2][14][13] = 3'b111;\
sp[2][14][14] = 3'b000;\
sp[2][14][15] = 3'b000;\
sp[2][15][0] = 3'b000;\
sp[2][15][1] = 3'b000;\
sp[2][15][2] = 3'b000;\
sp[2][15][3] = 3'b111;\
sp[2][15][4] = 3'b111;\
sp[2][15][5] = 3'b000;\
sp[2][15][6] = 3'b000;\
sp[2][15][7] = 3'b000;\
sp[2][15][8] = 3'b000;\
sp[2][15][9] = 3'b111;\
sp[2][15][10] = 3'b111;\
sp[2][15][11] = 3'b000;\
sp[2][15][12] = 3'b000;\
sp[2][15][13] = 3'b000;\
sp[2][15][14] = 3'b000;\
sp[2][15][15] = 3'b000;\
